// -----------------------------------------------------------------------------
// File        : packet_class.sv
// Author      : Varsha R (1BM23EC284)
// Created     : 2026-01-29
// Module      : packet_class
// Project     : SystemVerilog and Verification (23EC6PE2SV),
//               Faculty: Prof. Ajaykumar Devarapalli
// Description : a dummy module for the functionality.
// ----------------------------------------------------------------------------- 
module packet_class;
endmodule
